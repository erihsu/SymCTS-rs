module s1238_bench
(G2 , G546 , G535 , G8 , G547 , G5 , G537 , G530 , G45 , G549 , G0 , G12 , G548 , blif_clk_net , G539 , G3 , G13 , G552 , G6 , G542 , G4 , G10 , G9 , G1 , blif_reset_net , G11 , G550 , G532 , G551 , G7);
input G3;
input G2;
input G1;
input G0;
input blif_reset_net;
input blif_clk_net;
input G11;
input G10;
input G9;
input G8;
input G7;
input G6;
input G5;
input G4;
output G546;
output G542;
output G552;
output G551;
output G550;
output G549;
input G13;
input G12;
output G539;
output G45;
output G537;
output G535;
output G532;
output G530;
output G548;
output G547;
INV_X0P5B_A9TL40 U98 (.Y ( n668 ));
INV_X0P8M_A9TL40 U97 (.Y ( n667 ));
INV_X0P5B_A9TL40 U96 (.Y ( n666 ));
INV_X1M_A9TL40 U95 (.Y ( n665 ));
INV_X0P5B_A9TL40 U94 (.Y ( n664 ));
INV_X0P6M_A9TL40 U93 (.Y ( n663 ));
INV_X0P5B_A9TL40 U92 (.Y ( n662 ));
INV_X0P6M_A9TL40 U91 (.Y ( n661 ));
INV_X0P5B_A9TL40 U90 (.Y ( n660 ));
INV_X1B_A9TL40 U89 (.Y ( n659 ));
INV_X0P5B_A9TL40 U88 (.Y ( n658 ));
INV_X0P8M_A9TL40 U87 (.Y ( n657 ));
BUF_X1P2M_A9TL40 U86 (.Y ( n656 ));
INV_X0P5B_A9TL40 U85 (.Y ( n655 ));
INV_X0P7B_A9TL40 U84 (.Y ( n654 ));
INV_X0P5B_A9TL40 U83 (.Y ( n653 ));
INV_X0P7B_A9TL40 U82 (.A ( n653 ));
INV_X0P5B_A9TL40 U81 (.Y ( n651 ));
INV_X0P7B_A9TL40 U80 (.Y ( n650 ));
INV_X0P5B_A9TL40 U79 (.Y ( n649 ));
INV_X0P8M_A9TL40 U78 (.Y ( n648 ));
INV_X0P5B_A9TL40 U77 (.Y ( n647 ));
INV_X1M_A9TL40 U76 (.Y ( n646 ));
BUF_X1P2M_A9TL40 U75 (.Y ( n645 ));
INV_X0P5B_A9TL40 U74 (.Y ( n644 ));
INV_X0P7B_A9TL40 U73 (.A ( n644 ));
INV_X0P5B_A9TL40 U72 (.Y ( n642 ));
INV_X1B_A9TL40 U71 (.Y ( n641 ));
INV_X0P5B_A9TL40 U70 (.Y ( n640 ));
INV_X0P8M_A9TL40 U69 (.Y ( n639 ));
BUF_X1P2M_A9TL40 U68 (.Y ( n638 ));
INV_X0P5B_A9TL40 U67 (.Y ( n637 ));
INV_X0P8B_A9TL40 U66 (.Y ( n636 ));
INV_X0P5B_A9TL40 U65 (.Y ( n635 ));
INV_X0P6M_A9TL40 U64 (.Y ( n634 ));
INV_X0P5B_A9TL40 U63 (.Y ( n633 ));
INV_X0P6M_A9TL40 U62 (.Y ( n632 ));
INV_X0P5B_A9TL40 U61 (.Y ( n631 ));
INV_X0P8M_A9TL40 U60 (.Y ( n630 ));
INV_X0P5B_A9TL40 U22 (.Y ( n629 ));
INV_X0P5B_A9TL40 U59 (.Y ( n628 ));
INV_X1B_A9TL40 U58 (.Y ( n627 ));
INV_X0P5B_A9TL40 U57 (.Y ( n626 ));
INV_X1M_A9TL40 U56 (.Y ( n625 ));
INV_X0P5B_A9TL40 U55 (.Y ( n624 ));
INV_X1M_A9TL40 U54 (.Y ( n623 ));
INV_X0P5B_A9TL40 U53 (.Y ( n622 ));
INV_X1B_A9TL40 U52 (.Y ( n621 ));
INV_X0P5B_A9TL40 U51 (.Y ( n620 ));
INV_X1M_A9TL40 U50 (.Y ( n619 ));
INV_X0P5B_A9TL40 U49 (.Y ( n618 ));
INV_X1B_A9TL40 U48 (.Y ( n617 ));
INV_X0P5B_A9TL40 U47 (.Y ( n616 ));
INV_X0P7B_A9TL40 U46 (.Y ( n615 ));
BUF_X1P2M_A9TL40 U45 (.Y ( n614 ));
INV_X0P5B_A9TL40 U44 (.Y ( n613 ));
INV_X1B_A9TL40 U43 (.Y ( n612 ));
INV_X0P5B_A9TL40 U42 (.A ( n599 ));
INV_X1B_A9TL40 U41 (.Y ( n610 ));
INV_X0P5B_A9TL40 U40 (.Y ( n609 ));
INV_X0P8M_A9TL40 U39 (.Y ( n608 ));
INV_X0P5B_A9TL40 U38 (.Y ( n607 ));
INV_X0P7B_A9TL40 U37 (.Y ( n606 ));
INV_X0P5B_A9TL40 U36 (.Y ( n605 ));
INV_X0P8B_A9TL40 U35 (.Y ( n604 ));
INV_X0P5B_A9TL40 U24 (.Y ( n603 ));
INV_X1M_A9TL40 U23 (.Y ( n602 ));
INV_X1B_A9TL40 U4 (.Y ( n600 ));
BUF_X1P2M_A9TL40 U3 (.Y ( n599 ));
INV_X1B_A9TL40 U34 (.Y ( n598 ));
INV_X0P6B_A9TL40 U33 (.Y ( n597 ));
INV_X1B_A9TL40 U32 (.Y ( n596 ));
BUF_X1P2M_A9TL40 U31 (.Y ( n595 ));
INV_X0P8B_A9TL40 U30 (.Y ( n594 ));
BUF_X1P2M_A9TL40 U29 (.Y ( n593 ));
INV_X0P8B_A9TL40 U28 (.Y ( n592 ));
BUFH_X1M_A9TL40 U27 (.Y ( n591 ));
INV_X0P5B_A9TL40 U26 (.Y ( n590 ));
BUF_X1M_A9TL40 U25 (.Y ( n589 ));
INV_X0P8B_A9TL40 U21 (.Y ( n585 ));
BUF_X1M_A9TL40 U20 (.Y ( n584 ));
INV_X0P8B_A9TL40 U19 (.Y ( n583 ));
BUF_X1M_A9TL40 U18 (.Y ( n582 ));
INV_X0P8B_A9TL40 U17 (.Y ( n581 ));
BUFH_X1M_A9TL40 U16 (.Y ( n580 ));
INV_X0P5B_A9TL40 U15 (.Y ( n579 ));
BUFH_X1M_A9TL40 U14 (.Y ( n578 ));
INV_X0P5B_A9TL40 U13 (.Y ( n577 ));
BUF_X1M_A9TL40 U12 (.Y ( n576 ));
INV_X1B_A9TL40 U11 (.Y ( n575 ));
BUFH_X1M_A9TL40 U10 (.Y ( n574 ));
BUF_X1M_A9TL40 U9 (.Y ( n573 ));
INV_X0P8B_A9TL40 U8 (.Y ( n572 ));
BUFH_X1M_A9TL40 U7 (.Y ( n571 ));
INV_X1B_A9TL40 U6 (.Y ( n570 ));
BUF_X1M_A9TL40 U5 (.Y ( n569 ));
INV_X0P5B_A9TL40 U2 (.Y ( n566 ));
BUF_X1M_A9TL40 U1 (.A ( n625 ));
OAI31_X2M_A9TL40 U492 (.A1 ( n490 ) , .Y ( G530 ) , .A0 ( n589 ) , .A2 ( n495 ));
OAI211_X2M_A9TL40 U568 (.A0 ( n505 ) , .A1 ( n504 ) , .B0 ( n503 ) , .C0 ( n502 ));
AOI22_X1M_A9TL40 U423 (.Y ( n503 ) , .B1 ( n497 ) , .A1 ( n498 ) , .A0 ( n571 ));
INV_X1M_A9TL40 U302 (.Y ( n394 ));
AOI22_X1M_A9TL40 U352 (.Y ( n481 ) , .B1 ( n469 ) , .A1 ( n471 ) , .A0 ( n500 ));
NOR2_X0P5M_A9TL40 U331 (.Y ( n492 ) , .A ( n591 ));
AOI32_X1M_A9TL40 U459 (.A0 ( n441 ) , .A2 ( n312 ) , .Y ( n313 ) , .B0 ( n311 ) , .B1 ( n581 ));
NAND2_X3B_A9TL40 U533 (.Y ( n475 ) , .A ( n583 ));
INV_X0P5B_A9TL40 U332 (.Y ( n312 ));
NAND3_X0P5M_A9TL40 U441 (.Y ( n375 ) , .B ( n359 ) , .C ( n628 ));
NOR2_X0P5M_A9TL40 U421 (.Y ( n383 ) , .A ( n579 ));
NAND2_X0P5M_A9TL40 U471 (.Y ( n401 ) , .A ( n488 ));
NAND2_X0P5M_A9TL40 U412 (.Y ( n297 ) , .A ( n581 ));
INV_X0P5B_A9TL40 U321 (.Y ( n449 ));
INV_X0P5B_A9TL40 U557 (.Y ( n364 ));
INV_X0P5B_A9TL40 U320 (.Y ( n485 ));
NAND2_X0P5M_A9TL40 U481 (.Y ( n400 ) , .A ( n569 ));
NOR3_X0P5M_A9TL40 U411 (.Y ( n362 ) , .A ( n383 ) , .C ( n577 ));
NOR3_X0P5M_A9TL40 U417 (.Y ( n399 ) , .A ( n627 ) , .C ( n596 ));
OA1B2_X0P5M_A9TL40 U498 (.A0N ( n596 ) , .B1 ( n329 ) , .B0 ( n330 ));
NAND2_X0P5M_A9TL40 U538 (.Y ( n298 ) , .A ( n576 ));
NOR2_X0P5M_A9TL40 U489 (.Y ( n304 ) , .A ( n571 ));
NOR2_X0P5M_A9TL40 U488 (.Y ( n301 ) , .A ( n575 ));
NOR2_X0P5M_A9TL40 U543 (.Y ( n308 ) , .A ( n414 ));
NOR3_X0P5M_A9TL40 U496 (.Y ( n323 ) , .A ( n569 ) , .C ( n359 ));
NOR3_X0P5M_A9TL40 U497 (.Y ( n303 ) , .A ( n580 ) , .C ( n453 ));
NOR3_X0P5M_A9TL40 U303 (.Y ( n322 ) , .A ( n594 ) , .C ( n345 ));
INV_X0P5B_A9TL40 U528 (.Y ( G546 ));
INV_X0P5B_A9TL40 U299 (.Y ( n506 ));
NAND2_X0P5M_A9TL40 U361 (.Y ( G507 ) , .A ( n394 ));
NAND2_X0P5M_A9TL40 U544 (.Y ( G508 ) , .A ( n435 ));
INV_X0P5B_A9TL40 U545 (.Y ( n321 ));
NOR3_X1M_A9TL40 U546 (.Y ( n310 ) , .A ( n577 ) , .C ( n574 ));
NOR2_X0P7M_A9TL40 U540 (.Y ( n332 ) , .A ( n578 ));
NOR2_X1M_A9TL40 U526 (.Y ( n462 ) , .A ( n571 ));
NAND2_X0P5M_A9TL40 U535 (.Y ( n385 ) , .A ( n582 ));
NOR2_X1B_A9TL40 U328 (.Y ( n414 ) , .A ( n570 ));
NOR2_X0P5M_A9TL40 U530 (.Y ( n302 ) , .A ( n585 ));
NOR2_X0P5M_A9TL40 U527 (.Y ( n487 ) , .A ( n593 ));
AOI32_X0P7M_A9TL40 U548 (.A0 ( n315 ) , .A2 ( n314 ) , .Y ( n316 ) , .B0 ( n313 ) , .B1 ( n585 ));
INV_X0P5B_A9TL40 U468 (.Y ( n423 ));
INV_X0P5B_A9TL40 U479 (.Y ( n381 ));
AOI21_X0P7M_A9TL40 U549 (.Y ( n318 ) , .A1 ( n570 ) , .A0 ( n317 ));
OAI211_X0P5M_A9TL40 U551 (.A0 ( n380 ) , .A1 ( n321 ) , .B0 ( n320 ) , .C0 ( n360 ));
NOR2_X1B_A9TL40 U461 (.Y ( n353 ) , .A ( n495 ));
NAND2_X0P5M_A9TL40 U552 (.Y ( n345 ) , .A ( n328 ));
NOR3_X1M_A9TL40 U558 (.Y ( n428 ) , .A ( n627 ) , .C ( n359 ));
AOI22_X0P5M_A9TL40 U440 (.Y ( n407 ) , .B1 ( n462 ) , .A1 ( n493 ) , .A0 ( n592 ));
NAND2_X0P5M_A9TL40 U447 (.Y ( n369 ) , .A ( n345 ));
INV_X0P6M_A9TL40 U554 (.Y ( n482 ));
AND2_X0P5M_A9TL40 U356 (.A ( n395 ) , .Y ( n486 ));
NOR2_X0P5M_A9TL40 U362 (.Y ( n395 ) , .A ( n499 ));
NOR2_X1B_A9TL40 U438 (.Y ( n413 ) , .A ( n592 ));
NOR2_X1B_A9TL40 U367 (.Y ( n432 ) , .A ( n371 ));
NOR2_X0P5M_A9TL40 U297 (.Y ( n387 ) , .A ( n575 ));
NOR2_X0P5M_A9TL40 U439 (.Y ( n451 ) , .A ( n366 ));
INV_X0P5B_A9TL40 U559 (.Y ( n426 ));
NOR2_X0P5M_A9TL40 U360 (.Y ( n500 ) , .A ( n590 ));
AOI21_X0P5M_A9TL40 U433 (.Y ( n411 ) , .A1 ( n598 ) , .A0 ( n413 ));
NAND2_X0P7M_A9TL40 U437 (.Y ( n438 ) , .A ( n566 ));
AO21A1AI2_X0P5M_A9TL40 U567 (.Y ( n498 ) , .C0 ( n489 ) , .A1 ( n593 ) , .A0 ( n589 ));
AOI2XB1_X0P5M_A9TL40 U556 (.A0 ( n439 ) , .Y ( n476 ) , .B0 ( n565 ));
OA21A1OI2_X0P5M_A9TL40 U560 (.C0 ( n360 ) , .A0 ( n579 ) , .A1 ( n364 ) , .Y ( n422 ));
NOR2_X0P5M_A9TL40 U565 (.Y ( n470 ) , .A ( n595 ));
OAI211_X0P7M_A9TL40 U562 (.A0 ( G40 ) , .A1 ( n418 ) , .B0 ( n417 ) , .C0 ( n416 ));
OA21A1OI2_X0P5M_A9TL40 U566 (.C0 ( n470 ) , .A0 ( n486 ) , .A1 ( n433 ) , .Y ( n434 ));
NAND2_X0P5B_A9TL40 U476 (.Y ( n377 ) , .A ( n583 ));
NOR2_X1M_A9TL40 U477 (.Y ( n441 ) , .A ( n576 ));
AND4_X0P5M_A9TL40 U478 (.C ( n590 ) , .A ( n576 ) , .D ( n583 ) , .Y ( G511 ));
NAND2_X0P5B_A9TL40 U480 (.Y ( n406 ) , .A ( n596 ));
OA21_X0P5M_A9TL40 U482 (.A1 ( n577 ) , .B0 ( n383 ) , .Y ( n420 ));
NAND2_X0P5B_A9TL40 U483 (.Y ( n341 ) , .A ( n594 ));
OAI31_X1M_A9TL40 U485 (.A1 ( n330 ) , .Y ( n368 ) , .A0 ( n331 ) , .A2 ( n329 ));
NAND3_X0P5M_A9TL40 U486 (.Y ( n473 ) , .B ( n332 ) , .C ( n302 ));
NAND3_X0P5M_A9TL40 U490 (.Y ( n358 ) , .B ( n583 ) , .C ( n575 ));
OAI22_X0P5M_A9TL40 U491 (.Y ( G539 ) , .A0 ( n376 ) , .A1 ( n375 ) , .B1 ( n374 ));
OAI22_X0P5M_A9TL40 U493 (.Y ( G547 ) , .A0 ( n389 ) , .A1 ( n426 ) , .B1 ( n581 ));
NAND3_X0P5M_A9TL40 U494 (.Y ( n416 ) , .B ( n491 ) , .C ( n597 ));
NAND3_X0P5M_A9TL40 U495 (.Y ( n502 ) , .B ( n500 ) , .C ( n499 ));
OAI22_X0P5M_A9TL40 U499 (.Y ( n307 ) , .A0 ( n592 ) , .A1 ( n415 ) , .B1 ( n429 ));
OAI31_X0P5M_A9TL40 U500 (.A1 ( n574 ) , .Y ( n296 ) , .A0 ( n381 ) , .A2 ( n577 ));
AO21A1AI2_X0P5M_A9TL40 U501 (.Y ( G513 ) , .C0 ( n578 ) , .A1 ( n583 ) , .A0 ( n301 ));
AOI21_X0P5M_A9TL40 U502 (.Y ( G502 ) , .A1 ( n597 ) , .A0 ( n487 ));
NAND3_X0P5M_A9TL40 U503 (.Y ( n293 ) , .B ( n492 ) , .C ( n570 ));
OA21_X0P5M_A9TL40 U523 (.A1 ( n585 ) , .B0 ( n583 ) , .Y ( n287 ));
NAND3_X0P5M_A9TL40 U524 (.Y ( n490 ) , .B ( n428 ) , .C ( n596 ));
AO21A1AI2_X0P5M_A9TL40 U525 (.Y ( n291 ) , .C0 ( n591 ) , .A1 ( n570 ) , .A0 ( n595 ));
OAI21_X0P5M_A9TL40 U529 (.A1 ( n581 ) , .Y ( G510 ) , .B0 ( n297 ));
OAI22_X0P5M_A9TL40 U531 (.Y ( G504 ) , .A0 ( n576 ) , .A1 ( n585 ) , .B1 ( n583 ));
AOI22_X0P5M_A9TL40 U532 (.Y ( G512 ) , .B1 ( n594 ) , .A1 ( n598 ) , .A0 ( n593 ));
AOI21_X0P5M_A9TL40 U534 (.Y ( n295 ) , .A1 ( n449 ) , .A0 ( n383 ));
AOI22_X0P5M_A9TL40 U536 (.Y ( G515 ) , .B1 ( n385 ) , .A1 ( n296 ) , .A0 ( n584 ));
OAI211_X0P5M_A9TL40 U537 (.A0 ( n575 ) , .A1 ( n585 ) , .B0 ( n576 ) , .C0 ( n297 ));
AOI22_X0P5M_A9TL40 U539 (.Y ( n300 ) , .B1 ( n298 ) , .A1 ( n299 ) , .A0 ( n312 ));
NAND2XB_X0P5M_A9TL40 U541 (.Y ( G509 ) , .BN ( n304 ));
NAND2_X1M_A9TL40 U542 (.Y ( n495 ) , .A ( n571 ));
AOI211_X1M_A9TL40 U547 (.Y ( n311 ) , .C0 ( n310 ) , .A1 ( G31 ) , .A0 ( n578 ));
OAI211_X1M_A9TL40 U550 (.A0 ( n338 ) , .A1 ( n319 ) , .B0 ( G46 ) , .C0 ( n318 ));
NOR3_X1A_A9TL40 U553 (.Y ( n491 ) , .A ( n565 ) , .C ( n345 ));
NAND2_X0P5B_A9TL40 U555 (.Y ( n439 ) , .A ( n367 ));
OAI22_X0P5M_A9TL40 U561 (.Y ( G548 ) , .A0 ( n365 ) , .A1 ( n364 ) , .B1 ( n418 ));
OAI21_X0P5M_A9TL40 U563 (.A1 ( n585 ) , .Y ( n421 ) , .B0 ( n580 ));
NAND2_X0P5B_A9TL40 U564 (.Y ( n430 ) , .A ( n570 ));
NAND2_X0P5B_A9TL40 U383 (.Y ( n435 ) , .A ( n336 ));
NAND2XB_X0P5M_A9TL40 U384 (.Y ( n445 ) , .BN ( n454 ));
AOI211_X0P5M_A9TL40 U385 (.Y ( n505 ) , .C0 ( n483 ) , .A1 ( n572 ) , .A0 ( n485 ));
AO21A1AI2_X0P5M_A9TL40 U386 (.Y ( n288 ) , .C0 ( n589 ) , .A1 ( n597 ) , .A0 ( n341 ));
AOI21_X0P5M_A9TL40 U387 (.Y ( n327 ) , .A1 ( n390 ) , .A0 ( n598 ));
AOI22_X0P5M_A9TL40 U388 (.Y ( n342 ) , .B1 ( n575 ) , .A1 ( n336 ) , .A0 ( n467 ));
NAND2_X0P5B_A9TL40 U389 (.Y ( n472 ) , .A ( n572 ));
NOR3_X0P7M_A9TL40 U390 (.Y ( n467 ) , .A ( n572 ) , .C ( n390 ));
AOI21_X0P5M_A9TL40 U391 (.Y ( n365 ) , .A1 ( n363 ) , .A0 ( n584 ));
OAI22BB_X0P5M_A9TL40 U392 (.A1 ( n597 ) , .Y ( n393 ) , .B1N ( n487 ) , .B0N ( n571 ));
AOI21_X0P5M_A9TL40 U393 (.Y ( n389 ) , .A1 ( n380 ) , .A0 ( n381 ));
OAI31_X0P5M_A9TL40 U394 (.A1 ( n406 ) , .Y ( n335 ) , .A0 ( n571 ) , .A2 ( n334 ));
NOR3_X0P7M_A9TL40 U395 (.Y ( n330 ) , .A ( n574 ) , .C ( n594 ));
OAI22_X0P5M_A9TL40 U396 (.Y ( n348 ) , .A0 ( n591 ) , .A1 ( n347 ) , .B1 ( n410 ));
OAI22_X0P5M_A9TL40 U397 (.Y ( n402 ) , .A0 ( n488 ) , .A1 ( n495 ) , .B1 ( n401 ));
OAI211_X0P5M_A9TL40 U398 (.A0 ( n576 ) , .A1 ( n383 ) , .B0 ( G34 ) , .C0 ( n382 ));
NAND3_X0P7M_A9TL40 U399 (.Y ( n454 ) , .B ( n423 ) , .C ( n302 ));
OAI21_X0P5M_A9TL40 U400 (.A1 ( n378 ) , .Y ( n320 ) , .B0 ( n423 ));
NAND2_X0P5B_A9TL40 U401 (.Y ( n347 ) , .A ( n595 ));
OAI22_X0P5M_A9TL40 U402 (.Y ( n363 ) , .A0 ( n381 ) , .A1 ( n380 ) , .B1 ( n385 ));
AOI21_X0P5M_A9TL40 U403 (.Y ( n324 ) , .A1 ( n574 ) , .A0 ( n593 ));
NAND3B_X0P5M_A9TL40 U404 (.AN ( n338 ) , .B ( n572 ) , .Y ( n453 ));
AOI22_X0P5M_A9TL40 U405 (.Y ( n315 ) , .B1 ( n321 ) , .A1 ( n581 ) , .A0 ( n332 ));
AOI211_X0P5M_A9TL40 U406 (.Y ( n427 ) , .C0 ( n419 ) , .A1 ( n421 ) , .A0 ( n582 ));
AOI21_X0P5M_A9TL40 U407 (.Y ( n431 ) , .A1 ( n256 ) , .A0 ( n569 ));
NAND2_X0P5B_A9TL40 U408 (.Y ( n466 ) , .A ( n570 ));
OR2_X0P5M_A9TL40 U409 (.B ( n571 ) , .A ( n465 ));
NAND2_X0P5B_A9TL40 U410 (.Y ( n338 ) , .A ( n585 ));
NAND4_X0P7M_A9TL40 U413 (.B ( n337 ) , .D ( n570 ) , .Y ( n436 ) , .A ( n595 ));
NAND2_X0P5B_A9TL40 U414 (.Y ( n465 ) , .A ( n591 ));
NOR3_X0P7M_A9TL40 U415 (.Y ( n419 ) , .A ( n578 ) , .C ( n577 ));
NAND2_X0P5B_A9TL40 U416 (.Y ( n309 ) , .A ( n581 ));
NAND2_X0P5B_A9TL40 U418 (.Y ( n319 ) , .A ( n582 ));
NOR2_X0P7M_A9TL40 U419 (.Y ( n448 ) , .A ( n569 ));
AOI22_X0P5M_A9TL40 U420 (.Y ( n317 ) , .B1 ( n596 ) , .A1 ( n589 ) , .A0 ( n595 ));
OAI211_X0P7M_A9TL40 U422 (.A0 ( n427 ) , .A1 ( n426 ) , .B0 ( n425 ) , .C0 ( n424 ));
AOI31_X0P7M_A9TL40 U424 (.A0 ( n414 ) , .Y ( n417 ) , .A2 ( n495 ) , .B0 ( n412 ));
OAI211_X0P7M_A9TL40 U425 (.A0 ( G29 ) , .A1 ( n496 ) , .B0 ( n404 ) , .C0 ( n403 ));
OAI211_X0P5M_A9TL40 U426 (.A0 ( n398 ) , .A1 ( n504 ) , .B0 ( n397 ) , .C0 ( n396 ));
OAI211_X0P5M_A9TL40 U427 (.A0 ( G43 ) , .A1 ( n482 ) , .B0 ( n481 ) , .C0 ( n480 ));
AOI31_X0P7M_A9TL40 U428 (.A0 ( n431 ) , .Y ( n433 ) , .A2 ( n429 ) , .B0 ( n496 ));
OAI31_X0P7M_A9TL40 U429 (.A1 ( n496 ) , .Y ( n497 ) , .A0 ( n595 ) , .A2 ( n495 ));
OAI22_X0P7M_A9TL40 U430 (.Y ( n412 ) , .A0 ( n411 ) , .A1 ( n410 ) , .B1 ( n594 ));
AOI211_X0P7M_A9TL40 U431 (.Y ( n397 ) , .C0 ( n486 ) , .A1 ( n570 ) , .A0 ( n405 ));
OAI31_X0P5M_A9TL40 U432 (.A1 ( n478 ) , .Y ( n480 ) , .A0 ( n479 ) , .A2 ( n477 ));
NOR2XB_X0P7M_A9TL40 U434 (.A ( n437 ) , .BN ( G38 ));
OAI31_X0P7M_A9TL40 U435 (.A1 ( n418 ) , .Y ( n386 ) , .A0 ( n574 ) , .A2 ( n385 ));
OAI22_X0P7M_A9TL40 U436 (.Y ( n408 ) , .A0 ( n575 ) , .A1 ( n407 ) , .B1 ( n406 ));
INV_X0P6B_A9TL40 U442 (.Y ( n370 ));
NOR2XB_X0P5M_A9TL40 U443 (.A ( n628 ) , .BN ( n368 ));
NOR3_X2M_A9TL40 U444 (.Y ( n493 ) , .B ( n628 ) , .C ( n368 ));
OAI211_X0P7M_A9TL40 U445 (.A0 ( n342 ) , .A1 ( n341 ) , .B0 ( n340 ) , .C0 ( n445 ));
OAI31_X0P5M_A9TL40 U446 (.A1 ( n574 ) , .Y ( n290 ) , .A0 ( n582 ) , .A2 ( G30 ));
AO21A1AI2_X0P7M_A9TL40 U448 (.Y ( n366 ) , .C0 ( n591 ) , .A1 ( n335 ) , .A0 ( n337 ));
OAI31_X0P5M_A9TL40 U449 (.A1 ( n378 ) , .Y ( n356 ) , .A0 ( n351 ) , .A2 ( n377 ));
OA21A1OI2_X0P7M_A9TL40 U450 (.C0 ( n472 ) , .A0 ( n380 ) , .A1 ( n475 ) , .Y ( n344 ));
OAI21_X0P5M_A9TL40 U451 (.A1 ( n472 ) , .Y ( n447 ) , .B0 ( n445 ));
AOI31_X0P7M_A9TL40 U452 (.A0 ( n327 ) , .Y ( n331 ) , .A2 ( n391 ) , .B0 ( n592 ));
AOI211_X0P7M_A9TL40 U453 (.Y ( n355 ) , .C0 ( n474 ) , .A1 ( n354 ) , .A0 ( n454 ));
NAND2_X0P5B_A9TL40 U454 (.Y ( n351 ) , .A ( n592 ));
OAI22_X0P5M_A9TL40 U455 (.Y ( n456 ) , .A0 ( n597 ) , .A1 ( n454 ) , .B1 ( n453 ));
OAI211_X0P5M_A9TL40 U456 (.A0 ( n569 ) , .A1 ( n256 ) , .B0 ( n406 ) , .C0 ( n391 ));
AO21B_X0P5M_A9TL40 U457 (.A1 ( n467 ) , .Y ( n469 ) , .B0N ( n466 ));
AO21A1AI2_X0P5M_A9TL40 U458 (.Y ( n350 ) , .C0 ( n348 ) , .A1 ( n468 ) , .A0 ( n584 ));
OAI211_X0P5M_A9TL40 U460 (.A0 ( n569 ) , .A1 ( n465 ) , .B0 ( n464 ) , .C0 ( n463 ));
NAND2_X0P5B_A9TL40 U462 (.Y ( n391 ) , .A ( n571 ));
NAND2_X0P5B_A9TL40 U463 (.Y ( n382 ) , .A ( n578 ));
OAI211_X0P5M_A9TL40 U464 (.A0 ( n579 ) , .A1 ( n581 ) , .B0 ( n423 ) , .C0 ( G34 ));
INV_X0P6B_A9TL40 U465 (.Y ( n349 ));
OAI22_X0P5M_A9TL40 U466 (.Y ( n379 ) , .A0 ( n578 ) , .A1 ( n378 ) , .B1 ( n377 ));
AO21A1AI2_X0P5M_A9TL40 U467 (.Y ( n464 ) , .C0 ( n596 ) , .A1 ( n594 ) , .A0 ( n591 ));
OAI31_X0P5M_A9TL40 U469 (.A1 ( n596 ) , .Y ( n294 ) , .A0 ( n591 ) , .A2 ( n400 ));
NAND2_X0P7B_A9TL40 U470 (.Y ( n360 ) , .A ( n381 ));
NAND4XXXB_X1M_A9TL40 U472 (.A ( n578 ) , .Y ( n314 ) , .B ( n312 ) , .C ( n475 ));
AOI211_X0P7M_A9TL40 U473 (.Y ( n329 ) , .C0 ( n594 ) , .A1 ( n410 ) , .A0 ( n572 ));
NAND4_X0P5A_A9TL40 U474 (.B ( n332 ) , .D ( n581 ) , .Y ( n334 ) , .A ( n582 ));
OAI221_X0P5M_A9TL40 U475 (.B0 ( n594 ) , .A1 ( n598 ) , .A0 ( n593 ) , .Y ( n463 ) , .C0 ( n569 ));
INV_X0P6B_A9TL40 U290 (.Y ( n425 ));
AOI211_X0P5M_A9TL40 U291 (.Y ( G514 ) , .C0 ( n361 ) , .A1 ( n420 ) , .A0 ( G34 ));
INV_X0P6B_A9TL40 U292 (.Y ( n460 ));
AOI21_X0P5M_A9TL40 U293 (.Y ( n409 ) , .A1 ( n491 ) , .A0 ( n483 ));
INV_X0P7B_A9TL40 U294 (.Y ( n504 ));
INV_X0P6B_A9TL40 U295 (.Y ( n444 ));
INV_X0P7B_A9TL40 U296 (.Y ( n496 ));
OAI22_X0P5M_A9TL40 U298 (.Y ( n440 ) , .A0 ( n565 ) , .A1 ( n439 ) , .B1 ( n472 ));
INV_X0P6B_A9TL40 U300 (.Y ( n376 ));
OAI31_X1M_A9TL40 U301 (.A1 ( n436 ) , .Y ( n367 ) , .A0 ( n591 ) , .A2 ( n358 ));
NOR2_X0P7M_A9TL40 U304 (.Y ( n479 ) , .A ( n436 ));
INV_X0P6B_A9TL40 U305 (.Y ( n474 ));
INV_X0P7B_A9TL40 U306 (.Y ( n336 ));
NOR2_X0P5A_A9TL40 U307 (.Y ( n484 ) , .A ( n487 ));
INV_X0P6B_A9TL40 U308 (.Y ( n354 ));
NOR2_X0P7M_A9TL40 U309 (.Y ( n483 ) , .A ( n595 ));
NOR3_X0P5A_A9TL40 U310 (.Y ( n457 ) , .A ( n572 ) , .C ( n473 ));
OAI22_X0P5M_A9TL40 U311 (.Y ( n325 ) , .A0 ( n598 ) , .A1 ( n390 ) , .B1 ( n324 ));
INV_X0P7B_A9TL40 U312 (.Y ( n346 ));
AOI2XB1_X0P5M_A9TL40 U313 (.A0 ( n332 ) , .Y ( n446 ) , .B0 ( n468 ));
NOR2_X0P7M_A9TL40 U314 (.Y ( n352 ) , .A ( n475 ));
INV_X0P7B_A9TL40 U315 (.Y ( n339 ));
INV_X0P7B_A9TL40 U316 (.Y ( n499 ));
NAND4_X0P5A_A9TL40 U317 (.B ( n598 ) , .D ( G511 ) , .Y ( n333 ) , .A ( n578 ));
INV_X0P7B_A9TL40 U319 (.Y ( n390 ));
INV_X0P7B_A9TL40 U322 (.Y ( n326 ));
NOR2_X1B_A9TL40 U323 (.Y ( n488 ) , .A ( n570 ));
NAND2_X0P5B_A9TL40 U324 (.Y ( n415 ) , .A ( n574 ));
INV_X0P7B_A9TL40 U325 (.Y ( n410 ));
NOR3_X1M_A9TL40 U326 (.Y ( n468 ) , .A ( n582 ) , .C ( n309 ));
INV_X0P7B_A9TL40 U327 (.Y ( n380 ));
INV_X0P7B_A9TL40 U330 (.Y ( n378 ));
NOR2_X0P5A_A9TL40 U337 (.Y ( n337 ) , .A ( n585 ));
OR2_X0P7M_A9TL40 U343 (.B ( n596 ) , .A ( n572 ));
OAI211_X0P5M_A9TL40 U344 (.A0 ( G44 ) , .A1 ( n444 ) , .B0 ( n443 ) , .C0 ( n442 ));
OAI211_X0P5M_A9TL40 U345 (.A0 ( n461 ) , .A1 ( n460 ) , .B0 ( n459 ) , .C0 ( n458 ));
AOI22_X0P5M_A9TL40 U346 (.Y ( n403 ) , .B1 ( n402 ) , .A1 ( n486 ) , .A0 ( n595 ));
AOI22_X0P5M_A9TL40 U347 (.Y ( n443 ) , .B1 ( n450 ) , .A1 ( n479 ) , .A0 ( n476 ));
AOI31_X0P5M_A9TL40 U348 (.A0 ( n488 ) , .A2 ( n493 ) , .Y ( n489 ) , .B0 ( n486 ));
AOI22_X0P5M_A9TL40 U349 (.Y ( n459 ) , .B1 ( n449 ) , .A1 ( n451 ) , .A0 ( n452 ));
NAND2XB_X0P5M_A9TL40 U350 (.Y ( G518 ) , .BN ( n451 ));
OAI21_X0P5M_A9TL40 U351 (.A1 ( n468 ) , .Y ( n442 ) , .B0 ( n440 ));
OAI21_X0P5M_A9TL40 U353 (.A1 ( n456 ) , .Y ( n458 ) , .B0 ( n470 ));
AOI31_X0P5M_A9TL40 U354 (.A0 ( n582 ) , .A2 ( n387 ) , .Y ( n388 ) , .B0 ( n386 ));
OAI21_X0P5M_A9TL40 U355 (.A1 ( n405 ) , .Y ( n396 ) , .B0 ( n596 ));
NAND2_X0P5B_A9TL40 U357 (.Y ( n437 ) , .A ( n598 ));
AOI211_X0P5M_A9TL40 U358 (.Y ( n361 ) , .C0 ( n385 ) , .A1 ( n574 ) , .A0 ( n580 ));
AOI22_X0P5M_A9TL40 U359 (.Y ( n374 ) , .B1 ( n370 ) , .A1 ( n372 ) , .A0 ( n373 ));
INV_X0P6B_A9TL40 U363 (.Y ( n373 ));
AOI32_X0P5M_A9TL40 U364 (.A0 ( n589 ) , .A2 ( n323 ) , .Y ( G506 ) , .B0 ( n322 ) , .B1 ( n566 ));
AOI22_X0P5M_A9TL40 U365 (.Y ( n494 ) , .B1 ( G39 ) , .A1 ( n492 ) , .A0 ( n493 ));
AOI31_X0P5M_A9TL40 U366 (.A0 ( n593 ) , .A2 ( n291 ) , .Y ( n292 ) , .B0 ( n290 ));
NOR2_X1B_A9TL40 U368 (.Y ( n405 ) , .A ( n495 ));
AOI31_X1M_A9TL40 U369 (.A0 ( n584 ) , .A2 ( n594 ) , .Y ( n371 ) , .B0 ( n343 ));
AOI21_X0P5M_A9TL40 U370 (.Y ( n461 ) , .A1 ( n468 ) , .A0 ( n448 ));
AOI31_X0P5M_A9TL40 U371 (.A0 ( n491 ) , .A2 ( n400 ) , .Y ( n404 ) , .B0 ( n399 ));
AOI31_X0P5M_A9TL40 U372 (.A0 ( n593 ) , .A2 ( n356 ) , .Y ( n357 ) , .B0 ( n355 ));
AOI22_X0P5M_A9TL40 U373 (.Y ( n289 ) , .B1 ( n577 ) , .A1 ( n288 ) , .A0 ( n592 ));
AOI211_X0P5M_A9TL40 U374 (.Y ( G516 ) , .C0 ( n306 ) , .A1 ( n308 ) , .A0 ( n591 ));
AOI211_X0P5M_A9TL40 U375 (.Y ( n398 ) , .C0 ( n392 ) , .A1 ( n483 ) , .A0 ( n571 ));
NOR2_X0P5A_A9TL40 U376 (.Y ( n478 ) , .A ( n473 ));
OAI21_X0P5M_A9TL40 U377 (.A1 ( n495 ) , .Y ( G505 ) , .B0 ( n305 ));
NOR2_X0P7M_A9TL40 U378 (.Y ( n452 ) , .A ( n590 ));
NOR2_X0P5A_A9TL40 U379 (.Y ( n477 ) , .A ( n475 ));
AOI211_X0P5M_A9TL40 U380 (.Y ( G517 ) , .C0 ( n303 ) , .A1 ( n304 ) , .A0 ( n326 ));
AOI22_X0P5M_A9TL40 U381 (.Y ( n340 ) , .B1 ( n353 ) , .A1 ( G35 ) , .A0 ( n339 ));
AOI21_X0P5M_A9TL40 U382 (.Y ( n305 ) , .A1 ( n448 ) , .A0 ( n487 ));
DFFRPQ_X0P5M_A9TL40 G29_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G502 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G31_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G504 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G32_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G505 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G34_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G507 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G35_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G508 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G36_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G509 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G37_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G510 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G38_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G511 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G39_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G512 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G40_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G513 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G42_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G515 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G43_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G516 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G44_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G517 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G33_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G506 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G41_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G514 ) , .R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G45_reg (.CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .D ( G518 ) , .R ( n600 ));
DFFSQN_X0P5M_A9TL40 G46_reg (.D ( n506 ) , .CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .SN ( n629 ));
DFFSQN_X0P5M_A9TL40 G30_reg (.D ( n287 ) , .CK ( blif_clk_net_BUFH_X16M_A9TL40_0 ) , .SN ( n629 ));
INV_X1B_A9TL40 U289 (.Y ( n418 ));
BUFH_X16M_A9TL40 BUFH_X16M_A9TL40_0 (.Y ( blif_clk_net_BUFH_X16M_A9TL40_0 ));
endmodule
